`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
/*���ļ�Ϊ 32 λ 3 ѡ 1 MUX����ļ�
���룺
in_00��32 λ 00 �ڵ�����
in_01��32 λ 01 �ڵ�����
in_10��32 λ 10 �ڵ�����
sel��ѡ���ź�
�����
out ��MUX�����
*/
//////////////////////////////////////////////////////////////////////////////////


module MUX_32_3_1( 
in_00, in_01, in_10, sel, out
    );
    input[31:0] in_00, in_01, in_10;
    input[1:0] sel;
    output reg [31:0] out;
    
    always @ (*)
		begin
			case(sel)
				2'b00: out = in_00;
				2'b01: out = in_01;
				2'b10: out = in_10;
			endcase
		end
endmodule
