`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
/*���ļ�Ϊ 32 λ 2 ѡ 1 MUX�����ļ�
���룺

�����

*/
//////////////////////////////////////////////////////////////////////////////////


module SIM_MUX_32_2_1;
	reg sel;
	reg [31:0] x0;
	reg [31:0] x1;

	wire [31:0] y;

	MUX_2_1 mux_2_1_init(
		.in_0(x0), 
		.in_1(x1), 
		.sel(sel), 
		.out(y)
	);

	initial 
	   begin
	   
	   x0= 32'h0000FFF0; x1 = 32'h00000000; sel = 1'b0;
        #10 sel = 1'b0;x0 = 32'h00000000;
        #10 sel = 1'b0;x0 = 32'h00000000;
        #10 sel = 1'b1;x1 = 32'hFFFFFFFF;
        #10 sel = 1'b0;x1 = 32'h00F0F000;
        #10 $stop;

	   end
      
endmodule
