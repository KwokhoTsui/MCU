`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
/*���ļ�Ϊ 32 λ 3 ѡ 1 MUX�����ļ�
���룺

�����

*/
//////////////////////////////////////////////////////////////////////////////////


module SIM_MUX_32_3_1;
	reg [1:0]sel;
	reg [31:0] x00;
	reg [31:0] x01;
	reg [31:0] x10;

	wire [31:0] y;

	MUX_32_3_1 mux_3_1_init(
		.in_00(x00), 
		.in_01(x01), 
		.in_10(x10), 
		.sel(sel), 
		.out(y)
	);

	initial 
	   begin
	   
	   x00= 32'h0000FFF0; x01 = 32'h00000000; x10= 32'hFF00FFF0; sel = 2'b00;
        #10 sel = 2'b10;x10 = 32'h0F000000;
        #10 sel = 2'b00;x01 = 32'h00000000;
        #10 sel = 2'b10;x10 = 32'hFFFFFFFF;
        #10 sel = 2'b01;x00 = 32'h00F0F000;
        #10 $stop;

	   end
      
endmodule
