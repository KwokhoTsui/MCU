`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
/*���ļ���inst_mem�ķ����ļ�*/
//////////////////////////////////////////////////////////////////////////////////


module SIM_inst_mem;
    reg [31:0] A;
    wire [31:0] RD;
    
    inst_mem inst_mem_init(
    .A(A),
    .RD(RD)
    );
    
    initial 
	   begin
	   
	   A= 32'h00000000;
        #10 A = 32'h00000004;
        #10 A = 32'h0000000C;
        #10 A = 32'h00000010;
        #10 $stop;

	   end
	   
endmodule
